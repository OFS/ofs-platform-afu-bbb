//
// Placeholder file for the platform to copy in a pr_hssi_@group@_if.sv after
// the ofs_plat_if tree is generated. The placeholder causes the automatically
// generated platform_if_addenda files to load this file.
//
