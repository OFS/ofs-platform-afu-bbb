//
// Placeholder file for the platform to copy in a xCLASSx_xGROUPx_if.vh after
// the ofs_plat_if tree is generated. The placeholder causes the automatically
// generated platform_if_addenda files to put this directory on the include
// file list.
//
