//
// Copyright (c) 2020, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.

//
// Connect a pair of AXI stream interfaces with a skid buffer.
//

`include "ofs_plat_if.vh"

// Pass clock from slave to master
module ofs_plat_axi_stream_if_skid_slave_clk
   (
    ofs_plat_axi_stream_if.to_slave stream_slave,
    ofs_plat_axi_stream_if.to_master_clk stream_master
    );

    // synthesis translate_off
    `OFS_PLAT_AXI_STREAM_IF_CHECK_PARAMS_MATCH(stream_slave, stream_master)
    // synthesis translate_on

    assign stream_master.clk = stream_slave.clk;
    assign stream_master.reset_n = stream_slave.reset_n;
    // Debugging signal
    assign stream_master.instance_number = stream_slave.instance_number;

    ofs_plat_prim_ready_enable_skid
      #(
        .N_DATA_BITS(stream_master.T_PAYLOAD_WIDTH)
        )
      skid
       (
        .clk(stream_master.clk),
        .reset_n(stream_master.reset_n),

        .enable_from_src(stream_master.tvalid),
        .data_from_src(stream_master.t),
        .ready_to_src(stream_master.tready),

        .enable_to_dst(stream_slave.tvalid),
        .data_to_dst(stream_slave.t),
        .ready_from_dst(stream_slave.tready)
        );

endmodule // ofs_plat_axi_stream_if_skid_slave_clk


// Pass clock from master to slave
module ofs_plat_axi_stream_if_skid_master_clk
   (
    ofs_plat_axi_stream_if.to_slave_clk stream_slave,
    ofs_plat_axi_stream_if.to_master stream_master
    );

    // synthesis translate_off
    `OFS_PLAT_AXI_STREAM_IF_CHECK_PARAMS_MATCH(stream_slave, stream_master)
    // synthesis translate_on

    assign stream_slave.clk = stream_master.clk;
    assign stream_slave.reset_n = stream_master.reset_n;
    // Debugging signal
    assign stream_slave.instance_number = stream_master.instance_number;

    ofs_plat_prim_ready_enable_skid
      #(
        .N_DATA_BITS(stream_master.T_PAYLOAD_WIDTH)
        )
      skid
       (
        .clk(stream_master.clk),
        .reset_n(stream_master.reset_n),

        .enable_from_src(stream_master.tvalid),
        .data_from_src(stream_master.t),
        .ready_to_src(stream_master.tready),

        .enable_to_dst(stream_slave.tvalid),
        .data_to_dst(stream_slave.t),
        .ready_from_dst(stream_slave.tready)
        );

endmodule // ofs_plat_axi_stream_if_skid_master_clk
