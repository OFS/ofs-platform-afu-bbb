//
// Copyright (c) 2019, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.

`include "ofs_plat_if.vh"

//
// Map CCI-P MMIO requests to an Avalon memory channels. The AFU should supply
// the MMIO Avalon master.
//
// The MMIO data width must be a power of 2 between 64 and 512 bits. Addresses
// generated by the master here are to words (DATA_WIDTH). The data width of the
// word will affect the address size. Byteenable will indicate partial-word
// references.
//
// In CCI-P, the minimum addressable size is a DWORD.
//
module ofs_plat_map_ccip_as_avalon_mmio
  #(
    parameter MAX_OUTSTANDING_MMIO_RD_REQS = 64
    )
   (
    input  logic clk,
    input  logic reset,
    input  t_if_ccip_Rx sRx,
    output t_if_ccip_c2_Tx c2Tx,

    ofs_plat_avalon_mem_if.to_slave_clk mmio_to_afu
    );

    localparam DATA_WIDTH = mmio_to_afu.DATA_WIDTH_;
    typedef logic [DATA_WIDTH-1 : 0] t_mmio_data;

    localparam DATA_WIDTH_LEGAL = (DATA_WIDTH >= 64) && (DATA_WIDTH <= 512) &&
                                  (DATA_WIDTH == (2 ** $clog2(DATA_WIDTH)));
    // synthesis translate_off
    initial
    begin : error_proc
        if (! DATA_WIDTH_LEGAL)
            $fatal(2, "** ERROR ** %m: Data width (%0d) must be a power of 2 between 64 and 512.", DATA_WIDTH);
    end
    // synthesis translate_on

    assign mmio_to_afu.clk = clk;
    assign mmio_to_afu.reset = reset;

    // Index of the minimum addressable size (32 bit DWORD)
    localparam DWORD_IDX_BITS = $clog2(DATA_WIDTH / 32);
    typedef logic [DWORD_IDX_BITS-1 : 0] t_dword_idx;

    // Cast CCI-P c0 header into ReqMmioHdr
    t_ccip_c0_ReqMmioHdr mmio_in_hdr;
    assign mmio_in_hdr = t_ccip_c0_ReqMmioHdr'(sRx.c0.hdr);

    logic error;

    //
    // Send MMIO requests through a buffering FIFO in case the AFU's MMIO slave
    // asserts waitrequest.
    //
    logic req_in_fifo_notFull;
    logic mmio_is_wr;
    t_ccip_clData mmio_wr_data;
    t_ccip_c0_ReqMmioHdr mmio_hdr;
    logic mmio_req_deq;
    logic mmio_req_notEmpty;

    // Restructure incoming write data so that 32 and 64 bit writes are replicated
    // throughout, even in a 512 bit MMIO interface. Quartus will drop unused
    // replications.
    t_ccip_clData mmio_in_wr_data;
    always_comb
    begin
        if (mmio_in_hdr.length == 2'b00)
            // 32 bit write -- replicate 16 times
            mmio_in_wr_data = {16{sRx.c0.data[31:0]}};
        else if (mmio_in_hdr.length == 2'b01)
            // 64 bit write -- replicate 8 times
            mmio_in_wr_data = {8{sRx.c0.data[63:0]}};
        else
            // Full 512 bit write
            mmio_in_wr_data = sRx.c0.data[63:0];
    end

    ofs_plat_prim_fifo_bram
      #(
        // Simply push the whole data structures through the FIFO.
        // Quartus will remove the parts that wind up not being used.
        .N_DATA_BITS(1 + $bits(t_ccip_clData) + $bits(t_ccip_c0_ReqMmioHdr)),
        .N_ENTRIES(MAX_OUTSTANDING_MMIO_RD_REQS)
        )
      req_in_fifo
       (
        .clk,
        .reset,
        .enq_data({ sRx.c0.mmioWrValid, mmio_in_wr_data, mmio_in_hdr }),
        .enq_en((sRx.c0.mmioRdValid || sRx.c0.mmioWrValid) && ! error),
        .notFull(req_in_fifo_notFull),
        .almostFull(),
        .first({ mmio_is_wr, mmio_wr_data, mmio_hdr }),
        .deq_en(mmio_req_deq),
        .notEmpty(mmio_req_notEmpty)
        );

    //
    // Save tid for MMIO reads. It will be needed when generating the
    // response. Avalon slave responses will be returned in request order.
    //
    logic tid_in_fifo_notFull;
    t_ccip_tid mmio_tid;
    t_dword_idx dword_idx;

    ofs_plat_prim_fifo_bram
      #(
        .N_DATA_BITS($bits(t_dword_idx) + $bits(t_ccip_tid)),
        .N_ENTRIES(MAX_OUTSTANDING_MMIO_RD_REQS)
        )
      tid_in_fifo
       (
        .clk,
        .reset,
        .enq_data({ t_dword_idx'(mmio_in_hdr.address), mmio_in_hdr.tid }),
        .enq_en(sRx.c0.mmioRdValid && ! error),
        .notFull(tid_in_fifo_notFull),
        .almostFull(),
        .first({ dword_idx, mmio_tid }),
        .deq_en(mmio_to_afu.readdatavalid),
        // Must not be empty
        .notEmpty()
        );

    //
    // Ingress FIFO overflow check. Stop the FIFO if an overflow is detected.
    // This tends to be a far easier failure to debug than when an MMIO request
    // is dropped silently.
    //
    always_ff @(posedge clk)
    begin
        if (((sRx.c0.mmioRdValid || sRx.c0.mmioWrValid) && ! req_in_fifo_notFull) ||
            (sRx.c0.mmioRdValid && ! tid_in_fifo_notFull))
        begin
            error <= 1'b1;
        end

        if (reset)
        begin
            error <= !DATA_WIDTH_LEGAL;
        end
    end

    //
    // Generate requests to the MMIO slave.
    //
    assign mmio_to_afu.write = mmio_req_notEmpty && mmio_is_wr;
    assign mmio_to_afu.read = mmio_req_notEmpty && ! mmio_is_wr;
    assign mmio_to_afu.burstcount = 1;
    // Data has already been formatted properly for the mmio_to_afu word size.
    assign mmio_to_afu.writedata = t_mmio_data'(mmio_wr_data);

    // Drop low address bits. CCI-P's MMIO address space is to DWORDS. The Avalon
    // address space is the index of whatever the MMIO DATA_WIDTH is set to. The
    // low address bits will be reflected in byteenable.
    assign mmio_to_afu.address = mmio_hdr.address[$bits(t_ccip_mmioAddr)-1 : DWORD_IDX_BITS];

    typedef logic [(DATA_WIDTH/32)-1 : 0] t_dword_enable_mask;
    t_dword_enable_mask dword_enable_mask;

    typedef logic [(DATA_WIDTH/8)-1 : 0] t_byteenable;

    // Construct the byteenable mask based on the size and address of the request.
    always_comb
    begin
        // 512 bit access? This step leaves the mask all 1's if 512 bits and all 0's if not.
        dword_enable_mask = mmio_hdr.length[1] ? ~t_dword_enable_mask'(0) : t_dword_enable_mask'(0);

        // Now account for a 32 or 64 bit access. The mask here is one bit per 32 data
        // bits, since the minimum CCI-P reference encoding is 32 bits. This DWORD mask
        // will be expanded to the byteenable mask below.
        //
        // The index to dword_enable_mask is to 2 bit chunks of the mask, accounting for
        // aligned 64 bit requests. The low bit of t_dword_idx is forced to 0 to
        // guarantee alignment. Even for 32 bit requests, it selects the proper region
        // of dword_enable_mask. The value for the assignment is 2'b11 when masking a
        // 64 bit request and either 2'b10 or 2'b01 for 32 bit requests, depending on
        // which DWORD is being selected.
        //
        // This component is ORed into the mask to merge it with the 512 bit case above.
        dword_enable_mask[t_dword_idx'(mmio_hdr.address) & ~t_dword_idx'(1) +: 2] |=
            (mmio_hdr.length[0] ? 2'b11 : (mmio_hdr.address[0] ? 2'b10 : 2'b01));

        // Expand the dword_enable_mask to a byte enable mask
        for (int i = 0; i < $bits(t_dword_enable_mask); i = i + 1)
        begin : be
            mmio_to_afu.byteenable[4*i +: 4] = {4{dword_enable_mask[i]}};
        end
    end

    // Forward read responses back to CCI-P.
    always_ff @(posedge clk)
    begin
        c2Tx.mmioRdValid <= mmio_to_afu.readdatavalid;
        c2Tx.hdr.tid <= mmio_tid;

        c2Tx.data <= mmio_to_afu.readdata;
        if (dword_idx[0])
        begin
            c2Tx.data[31:0] <= mmio_to_afu.readdata[63:32];
        end

        if (reset)
        begin
            c2Tx.mmioRdValid <= 1'b0;
        end
    end


    //
    // Generate requests to the 512 bit slave.
    //
    // Convert to 512 bit words (from 32 bit words)
    //assign mmio512_wr_to_afu.address = mmio_hdr.address[$bits(t_ccip_mmioAddr)-1 : 4];


    //
    // Consume requests once they are accepted by the Avalon slave.
    //
    assign mmio_req_deq = ! mmio_to_afu.waitrequest && mmio_req_notEmpty;

endmodule // ofs_plat_map_ccip_as_avalon_mmio
