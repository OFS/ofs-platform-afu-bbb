// Copyright (C) 2022 Intel Corporation
// SPDX-License-Identifier: MIT

//
// Included for compatibility with legacy platform support. Modules may use
// either the OFS or the OPAE SDK platform interface.
//

`ifndef __PLATFORM_IF_VH__
`define __PLATFORM_IF_VH__

`include "ofs_plat_if.vh"

`endif
